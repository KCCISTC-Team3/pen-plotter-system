`timescale 1ns / 1ps

module Pixel_Clk_Gen (
    input  logic clk,
    input  logic reset,
    output logic pclk
);
    logic [2:0] p_counter;

    always_ff @(posedge clk, posedge reset) begin
        if (reset) begin
            p_counter <= 0;
        end else begin
            if (p_counter == 4) begin
                p_counter <= 0;
                pclk      <= 1'b1;
            end else begin
                p_counter <= p_counter + 1;
                pclk      <= 1'b0;
            end
        end
    end
endmodule
