module top_uart_tx_logic (
    input  logic       clk,
    input  logic       reset,
    input  logic       canny_de,
    input  logic [7:0] canny_data,
    output logic       tx

);

    logic                    we;
    logic [             7:0] wData;
    logic [$clog2(5100)-1:0] wAddr;
    logic                    frame_tick;
    logic                    tx_fifo_full;
    logic [             7:0] tx_data;

    pixel_8_fsm U_PIXEL_8_FSM (
        .clk       (clk),
        .reset     (reset),
        .canny_de  (canny_de),
        .canny_data(canny_data),
        .we        (we),
        .wData     (wData),
        .wAddr     (wAddr),
        .frame_tick(frame_tick)
    );

    tx_ram U_TX_RAM (
        .clk       (clk),
        .reset     (reset),
        .we        (we),
        .wData     (wData),
        .wAddr     (wAddr),
        .frame_tick(frame_tick),
        .re        (frame_done && ~tx_fifo_full),
        .rData     (tx_data),
        .frame_done(frame_done)
    );

    uart_tx_fifo U_UART_TX_FIFO (
        .clk         (clk),
        .reset       (reset),
        .tx_data     (tx_data),
        .push        (frame_done && ~tx_fifo_full),
        .tx          (tx),
        .tx_fifo_full(tx_fifo_full)
    );

endmodule

