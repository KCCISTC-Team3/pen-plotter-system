`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2026/01/06 11:34:48
// Design Name: 
// Module Name: data_assembly_fsm
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module data_assembly_fsm(
    input empty,
    input [7:0]pop_data,
    output [23:0]rgb_data,
    output       rgb_done,
    output       start,
    output       stop
    );
    
    
    
endmodule
